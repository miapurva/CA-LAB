module multiplier(x,y,o);

input [31:0]x,y;
//input clk;
output [64:0]o;
output [63:0]s1,s2,s3,s4,s5,s6,s7,s8,s9,s10,s11,s12,s13,s14,s15,s16,s17,s18,s19,s20,s21,s22,s23,s24,s25,s26,s27,s28,s29;
wire [63:0]p[31:0];
wire cout1,cout2;
output [63:0]c1,c2,c3,c4,c5,c6,c7,c8,c9,c10,c11,c12,c13,c14,c15,c16,c17,c18,c19,c20,c21,c22,c23,c24,c25,c26,c27,c28,c29,c30,s30;
//level 1
//assign p[0][31:0]=x[31:0] & y[0];
assign p[0][0] = x[0]&y[0];
assign p[0][1] = x[1]&y[0];
assign p[0][2] = x[2]&y[0];
assign p[0][3] = x[3]&y[0];
assign p[0][4] = x[4]&y[0];
assign p[0][5] = x[5]&y[0];
assign p[0][6] = x[6]&y[0];
assign p[0][7] = x[7]&y[0];
assign p[0][8] = x[8]&y[0];
assign p[0][9] = x[9]&y[0];
assign p[0][10] = x[10]&y[0];
assign p[0][11] = x[11]&y[0];
assign p[0][12] = x[12]&y[0];
assign p[0][13] = x[13]&y[0];
assign p[0][14] = x[14]&y[0];
assign p[0][15] = x[15]&y[0];
assign p[0][16] = x[16]&y[0];
assign p[0][17] = x[17]&y[0];
assign p[0][18] = x[18]&y[0];
assign p[0][19] = x[19]&y[0];
assign p[0][20] = x[20]&y[0];
assign p[0][21] = x[21]&y[0];
assign p[0][22] = x[22]&y[0];
assign p[0][23] = x[23]&y[0];
assign p[0][24] = x[24]&y[0];
assign p[0][25] = x[25]&y[0];
assign p[0][26] = x[26]&y[0];
assign p[0][27] = x[27]&y[0];
assign p[0][28] = x[28]&y[0];
assign p[0][29] = x[29]&y[0];
assign p[0][30] = x[30]&y[0];
assign p[0][31] = x[31]&y[0];
assign p[0][63:32]=1'b0;

//level 2
assign p[1][0] = 1'b0;
assign p[1][1] = x[0]&y[1];
assign p[1][2] = x[1]&y[1];
assign p[1][3] = x[2]&y[1];
assign p[1][4] = x[3]&y[1];
assign p[1][5] = x[4]&y[1];
assign p[1][6] = x[5]&y[1];
assign p[1][7] = x[6]&y[1];
assign p[1][8] = x[7]&y[1];
assign p[1][9] = x[8]&y[1];
assign p[1][10] = x[9]&y[1];
assign p[1][11] = x[10]&y[1];
assign p[1][12] = x[11]&y[1];
assign p[1][13] = x[12]&y[1];
assign p[1][14] = x[13]&y[1];
assign p[1][15] = x[14]&y[1];
assign p[1][16] = x[15]&y[1];
assign p[1][17] = x[16]&y[1];
assign p[1][18] = x[17]&y[1];
assign p[1][19] = x[18]&y[1];
assign p[1][20] = x[19]&y[1];
assign p[1][21] = x[20]&y[1];
assign p[1][22] = x[21]&y[1];
assign p[1][23] = x[22]&y[1];
assign p[1][24] = x[23]&y[1];
assign p[1][25] = x[24]&y[1];
assign p[1][26] = x[25]&y[1];
assign p[1][27] = x[26]&y[1];
assign p[1][28] = x[27]&y[1];
assign p[1][29] = x[28]&y[1];
assign p[1][30] = x[29]&y[1];
assign p[1][31] = x[30]&y[1];
assign p[1][32] = x[31]&y[1];
assign p[1][63:33]=1'b0;

//level3
assign p[2][1:0]=1'b0;
assign p[2][2]=x[0] & y[2];
assign p[2][3] = x[1]&y[2];
assign p[2][4] = x[2]&y[2];
assign p[2][5] = x[3]&y[2];
assign p[2][6] = x[4]&y[2];
assign p[2][7] = x[5]&y[2];
assign p[2][8] = x[6]&y[2];
assign p[2][9] = x[7]&y[2];
assign p[2][10] = x[8]&y[2];
assign p[2][11] = x[9]&y[2];
assign p[2][12] = x[10]&y[2];
assign p[2][13] = x[11]&y[2];
assign p[2][14] = x[12]&y[2];
assign p[2][15] = x[13]&y[2];
assign p[2][16] = x[14]&y[2];
assign p[2][17] = x[15]&y[2];
assign p[2][18] = x[16]&y[2];
assign p[2][19] = x[17]&y[2];
assign p[2][20] = x[18]&y[2];
assign p[2][21] = x[19]&y[2];
assign p[2][22] = x[20]&y[2];
assign p[2][23] = x[21]&y[2];
assign p[2][24] = x[22]&y[2];
assign p[2][25] = x[23]&y[2];
assign p[2][26] = x[24]&y[2];
assign p[2][27] = x[25]&y[2];
assign p[2][28] = x[26]&y[2];
assign p[2][29] = x[27]&y[2];
assign p[2][30] = x[28]&y[2];
assign p[2][31] = x[29]&y[2];
assign p[2][32] = x[30]&y[2];
assign p[2][33] = x[31]&y[2];
assign p[2][63:34]=1'b0;

//level4
assign p[3][2:0]=1'b0;
assign p[3][3]=x[0] & y[3];
assign p[3][4] = x[1]&y[3];
assign p[3][5] = x[2]&y[3];
assign p[3][6] = x[3]&y[3];
assign p[3][7] = x[4]&y[3];
assign p[3][8] = x[5]&y[3];
assign p[3][9] = x[6]&y[3];
assign p[3][10] = x[7]&y[3];
assign p[3][11] = x[8]&y[3];
assign p[3][12] = x[9]&y[3];
assign p[3][13] = x[10]&y[3];
assign p[3][14] = x[11]&y[3];
assign p[3][15] = x[12]&y[3];
assign p[3][16] = x[13]&y[3];
assign p[3][17] = x[14]&y[3];
assign p[3][18] = x[15]&y[3];
assign p[3][19] = x[16]&y[3];
assign p[3][20] = x[17]&y[3];
assign p[3][21] = x[18]&y[3];
assign p[3][22] = x[19]&y[3];
assign p[3][23] = x[20]&y[3];
assign p[3][24] = x[21]&y[3];
assign p[3][25] = x[22]&y[3];
assign p[3][26] = x[23]&y[3];
assign p[3][27] = x[24]&y[3];
assign p[3][28] = x[25]&y[3];
assign p[3][29] = x[26]&y[3];
assign p[3][30] = x[27]&y[3];
assign p[3][31] = x[28]&y[3];
assign p[3][32] = x[29]&y[3];
assign p[3][33] = x[30]&y[3];
assign p[3][34] = x[31]&y[3];
assign p[3][63:35]=1'b0;

//level5
assign p[4][3:0]=1'b0;
assign p[4][4]=x[0] & y[4];
assign p[4][5]=x[1] & y[4];
assign p[4][6] = x[2]&y[4];
assign p[4][7] = x[3]&y[4];
assign p[4][8] = x[4]&y[4];
assign p[4][9] = x[5]&y[4];
assign p[4][10] = x[6]&y[4];
assign p[4][11] = x[7]&y[4];
assign p[4][12] = x[8]&y[4];
assign p[4][13] = x[9]&y[4];
assign p[4][14] = x[10]&y[4];
assign p[4][15] = x[11]&y[4];
assign p[4][16] = x[12]&y[4];
assign p[4][17] = x[13]&y[4];
assign p[4][18] = x[14]&y[4];
assign p[4][19] = x[15]&y[4];
assign p[4][20] = x[16]&y[4];
assign p[4][21] = x[17]&y[4];
assign p[4][22] = x[18]&y[4];
assign p[4][23] = x[19]&y[4];
assign p[4][24] = x[20]&y[4];
assign p[4][25] = x[21]&y[4];
assign p[4][26] = x[22]&y[4];
assign p[4][27] = x[23]&y[4];
assign p[4][28] = x[24]&y[4];
assign p[4][29] = x[25]&y[4];
assign p[4][30] = x[26]&y[4];
assign p[4][31] = x[27]&y[4];
assign p[4][32] = x[28]&y[4];
assign p[4][33] = x[29]&y[4];
assign p[4][34] = x[30]&y[4];
assign p[4][35] = x[31]&y[4];
assign p[4][63:36]=1'b0;

//level6
assign p[5][4:0]=1'b0;
assign p[5][5] = x[0] & y[5];
assign p[5][6] = x[1]&y[5];
assign p[5][7] = x[2]&y[5];
assign p[5][8] = x[3]&y[5];
assign p[5][9] = x[4]&y[5];
assign p[5][10] = x[5]&y[5];
assign p[5][11] = x[6]&y[5];
assign p[5][12] = x[7]&y[5];
assign p[5][13] = x[8]&y[5];
assign p[5][14] = x[9]&y[5];
assign p[5][15] = x[10]&y[5];
assign p[5][16] = x[11]&y[5];
assign p[5][17] = x[12]&y[5];
assign p[5][18] = x[13]&y[5];
assign p[5][19] = x[14]&y[5];
assign p[5][20] = x[15]&y[5];
assign p[5][21] = x[16]&y[5];
assign p[5][22] = x[17]&y[5];
assign p[5][23] = x[18]&y[5];
assign p[5][24] = x[19]&y[5];
assign p[5][25] = x[20]&y[5];
assign p[5][26] = x[21]&y[5];
assign p[5][27] = x[22]&y[5];
assign p[5][28] = x[23]&y[5];
assign p[5][29] = x[24]&y[5];
assign p[5][30] = x[25]&y[5];
assign p[5][31] = x[26]&y[5];
assign p[5][32] = x[27]&y[5];
assign p[5][33] = x[28]&y[5];
assign p[5][34] = x[29]&y[5];
assign p[5][35] = x[30]&y[5];
assign p[5][36] = x[31]&y[5];
assign p[5][63:37]=1'b0;

//level7
assign p[6][5:0]=1'b0;
assign p[6][6]= x[0] & y[6];
assign p[6][7] = x[1]&y[6];
assign p[6][8] = x[2]&y[6];
assign p[6][9] = x[3]&y[6];
assign p[6][10] = x[4]&y[6];
assign p[6][11] = x[5]&y[6];
assign p[6][12] = x[6]&y[6];
assign p[6][13] = x[7]&y[6];
assign p[6][14] = x[8]&y[6];
assign p[6][15] = x[9]&y[6];
assign p[6][16] = x[10]&y[6];
assign p[6][17] = x[11]&y[6];
assign p[6][18] = x[12]&y[6];
assign p[6][19] = x[13]&y[6];
assign p[6][20] = x[14]&y[6];
assign p[6][21] = x[15]&y[6];
assign p[6][22] = x[16]&y[6];
assign p[6][23] = x[17]&y[6];
assign p[6][24] = x[18]&y[6];
assign p[6][25] = x[19]&y[6];
assign p[6][26] = x[20]&y[6];
assign p[6][27] = x[21]&y[6];
assign p[6][28] = x[22]&y[6];
assign p[6][29] = x[23]&y[6];
assign p[6][30] = x[24]&y[6];
assign p[6][31] = x[25]&y[6];
assign p[6][32] = x[26]&y[6];
assign p[6][33] = x[27]&y[6];
assign p[6][34] = x[28]&y[6];
assign p[6][35] = x[29]&y[6];
assign p[6][36] = x[30]&y[6];
assign p[6][37] = x[31]&y[6];
assign p[6][63:38]=1'b0;

//level8
assign p[7][6:0]=1'b0;
assign p[7][7]= x[0] & y[7];
assign p[7][8] = x[1]&y[7];
assign p[7][9] = x[2]&y[7];
assign p[7][10] = x[3]&y[7];
assign p[7][11] = x[4]&y[7];
assign p[7][12] = x[5]&y[7];
assign p[7][13] = x[6]&y[7];
assign p[7][14] = x[7]&y[7];
assign p[7][15] = x[8]&y[7];
assign p[7][16] = x[9]&y[7];
assign p[7][17] = x[10]&y[7];
assign p[7][18] = x[11]&y[7];
assign p[7][19] = x[12]&y[7];
assign p[7][20] = x[13]&y[7];
assign p[7][21] = x[14]&y[7];
assign p[7][22] = x[15]&y[7];
assign p[7][23] = x[16]&y[7];
assign p[7][24] = x[17]&y[7];
assign p[7][25] = x[18]&y[7];
assign p[7][26] = x[19]&y[7];
assign p[7][27] = x[20]&y[7];
assign p[7][28] = x[21]&y[7];
assign p[7][29] = x[22]&y[7];
assign p[7][30] = x[23]&y[7];
assign p[7][31] = x[24]&y[7];
assign p[7][32] = x[25]&y[7];
assign p[7][33] = x[26]&y[7];
assign p[7][34] = x[27]&y[7];
assign p[7][35] = x[28]&y[7];
assign p[7][36] = x[29]&y[7];
assign p[7][37] = x[30]&y[7];
assign p[7][38] = x[31]&y[7];
assign p[7][63:39]= 1'b0;

//level9
assign p[8][7:0]= 1'b0;
assign p[8][8] = x[0] & y[8];
assign p[8][9] = x[1]&y[8];
assign p[8][10] = x[2]&y[8];
assign p[8][11] = x[3]&y[8];
assign p[8][12] = x[4]&y[8];
assign p[8][13] = x[5]&y[8];
assign p[8][14] = x[6]&y[8];
assign p[8][15] = x[7]&y[8];
assign p[8][16] = x[8]&y[8];
assign p[8][17] = x[9]&y[8];
assign p[8][18] = x[10]&y[8];
assign p[8][19] = x[11]&y[8];
assign p[8][20] = x[12]&y[8];
assign p[8][21] = x[13]&y[8];
assign p[8][22] = x[14]&y[8];
assign p[8][23] = x[15]&y[8];
assign p[8][24] = x[16]&y[8];
assign p[8][25] = x[17]&y[8];
assign p[8][26] = x[18]&y[8];
assign p[8][27] = x[19]&y[8];
assign p[8][28] = x[20]&y[8];
assign p[8][29] = x[21]&y[8];
assign p[8][30] = x[22]&y[8];
assign p[8][31] = x[23]&y[8];
assign p[8][32] = x[24]&y[8];
assign p[8][33] = x[25]&y[8];
assign p[8][34] = x[26]&y[8];
assign p[8][35] = x[27]&y[8];
assign p[8][36] = x[28]&y[8];
assign p[8][37] = x[29]&y[8];
assign p[8][38] = x[30]&y[8];
assign p[8][39] = x[31]&y[8];
assign p[8][63:40] =1'b0;

//level 10
assign p[9][8:0]= 1'b0;
assign p[9][9] = x[0] & y[9];
assign p[9][10] = x[1]&y[9];
assign p[9][11] = x[2]&y[9];
assign p[9][12] = x[3]&y[9];
assign p[9][13] = x[4]&y[9];
assign p[9][14] = x[5]&y[9];
assign p[9][15] = x[6]&y[9];
assign p[9][16] = x[7]&y[9];
assign p[9][17] = x[8]&y[9];
assign p[9][18] = x[9]&y[9];
assign p[9][19] = x[10]&y[9];
assign p[9][20] = x[11]&y[9];
assign p[9][21] = x[12]&y[9];
assign p[9][22] = x[13]&y[9];
assign p[9][23] = x[14]&y[9];
assign p[9][24] = x[15]&y[9];
assign p[9][25] = x[16]&y[9];
assign p[9][26] = x[17]&y[9];
assign p[9][27] = x[18]&y[9];
assign p[9][28] = x[19]&y[9];
assign p[9][29] = x[20]&y[9];
assign p[9][30] = x[21]&y[9];
assign p[9][31] = x[22]&y[9];
assign p[9][32] = x[23]&y[9];
assign p[9][33] = x[24]&y[9];
assign p[9][34] = x[25]&y[9];
assign p[9][35] = x[26]&y[9];
assign p[9][36] = x[27]&y[9];
assign p[9][37] = x[28]&y[9];
assign p[9][38] = x[29]&y[9];
assign p[9][39] = x[30]&y[9];
assign p[9][40] = x[31]&y[9];
assign p[9][63:41] =1'b0;

//level 11
assign p[10][9:0]= 1'b0;
assign p[10][10] = x[0] & y[10];
assign p[10][11] = x[1]&y[10];
assign p[10][12] = x[2]&y[10];
assign p[10][13] = x[3]&y[10];
assign p[10][14] = x[4]&y[10];
assign p[10][15] = x[5]&y[10];
assign p[10][16] = x[6]&y[10];
assign p[10][17] = x[7]&y[10];
assign p[10][18] = x[8]&y[10];
assign p[10][19] = x[9]&y[10];
assign p[10][20] = x[10]&y[10];
assign p[10][21] = x[11]&y[10];
assign p[10][22] = x[12]&y[10];
assign p[10][23] = x[13]&y[10];
assign p[10][24] = x[14]&y[10];
assign p[10][25] = x[15]&y[10];
assign p[10][26] = x[16]&y[10];
assign p[10][27] = x[17]&y[10];
assign p[10][28] = x[18]&y[10];
assign p[10][29] = x[19]&y[10];
assign p[10][30] = x[20]&y[10];
assign p[10][31] = x[21]&y[10];
assign p[10][32] = x[22]&y[10];
assign p[10][33] = x[23]&y[10];
assign p[10][34] = x[24]&y[10];
assign p[10][35] = x[25]&y[10];
assign p[10][36] = x[26]&y[10];
assign p[10][37] = x[27]&y[10];
assign p[10][38] = x[28]&y[10];
assign p[10][39] = x[29]&y[10];
assign p[10][40] = x[30]&y[10];
assign p[10][41] = x[31]&y[10];
assign p[10][63:42] =1'b0;

//level 12
assign p[11][10:0]= 1'b0;
assign p[11][11] = x[0] & y[11];
assign p[11][12] = x[1]&y[11];
assign p[11][13] = x[2]&y[11];
assign p[11][14] = x[3]&y[11];
assign p[11][15] = x[4]&y[11];
assign p[11][16] = x[5]&y[11];
assign p[11][17] = x[6]&y[11];
assign p[11][18] = x[7]&y[11];
assign p[11][19] = x[8]&y[11];
assign p[11][20] = x[9]&y[11];
assign p[11][21] = x[10]&y[11];
assign p[11][22] = x[11]&y[11];
assign p[11][23] = x[12]&y[11];
assign p[11][24] = x[13]&y[11];
assign p[11][25] = x[14]&y[11];
assign p[11][26] = x[15]&y[11];
assign p[11][27] = x[16]&y[11];
assign p[11][28] = x[17]&y[11];
assign p[11][29] = x[18]&y[11];
assign p[11][30] = x[19]&y[11];
assign p[11][31] = x[20]&y[11];
assign p[11][32] = x[21]&y[11];
assign p[11][33] = x[22]&y[11];
assign p[11][34] = x[23]&y[11];
assign p[11][35] = x[24]&y[11];
assign p[11][36] = x[25]&y[11];
assign p[11][37] = x[26]&y[11];
assign p[11][38] = x[27]&y[11];
assign p[11][39] = x[28]&y[11];
assign p[11][40] = x[29]&y[11];
assign p[11][41] = x[30]&y[11];
assign p[11][42] = x[31]&y[11];
assign p[11][63:43] =1'b0;

//level 13
assign p[12][11:0]= 1'b0;
assign p[12][12] = x[0] & y[12];
assign p[12][13] = x[1]&y[12];
assign p[12][14] = x[2]&y[12];
assign p[12][15] = x[3]&y[12];
assign p[12][16] = x[4]&y[12];
assign p[12][17] = x[5]&y[12];
assign p[12][18] = x[6]&y[12];
assign p[12][19] = x[7]&y[12];
assign p[12][20] = x[8]&y[12];
assign p[12][21] = x[9]&y[12];
assign p[12][22] = x[10]&y[12];
assign p[12][23] = x[11]&y[12];
assign p[12][24] = x[12]&y[12];
assign p[12][25] = x[13]&y[12];
assign p[12][26] = x[14]&y[12];
assign p[12][27] = x[15]&y[12];
assign p[12][28] = x[16]&y[12];
assign p[12][29] = x[17]&y[12];
assign p[12][30] = x[18]&y[12];
assign p[12][31] = x[19]&y[12];
assign p[12][32] = x[20]&y[12];
assign p[12][33] = x[21]&y[12];
assign p[12][34] = x[22]&y[12];
assign p[12][35] = x[23]&y[12];
assign p[12][36] = x[24]&y[12];
assign p[12][37] = x[25]&y[12];
assign p[12][38] = x[26]&y[12];
assign p[12][39] = x[27]&y[12];
assign p[12][40] = x[28]&y[12];
assign p[12][41] = x[29]&y[12];
assign p[12][42] = x[30]&y[12];
assign p[12][43] = x[31]&y[12];
assign p[12][63:44] =1'b0;

//level 14
assign p[13][12:0]= 1'b0;
assign p[13][13] = x[0] & y[13];
assign p[13][14] = x[1]&y[13];
assign p[13][15] = x[2]&y[13];
assign p[13][16] = x[3]&y[13];
assign p[13][17] = x[4]&y[13];
assign p[13][18] = x[5]&y[13];
assign p[13][19] = x[6]&y[13];
assign p[13][20] = x[7]&y[13];
assign p[13][21] = x[8]&y[13];
assign p[13][22] = x[9]&y[13];
assign p[13][23] = x[10]&y[13];
assign p[13][24] = x[11]&y[13];
assign p[13][25] = x[12]&y[13];
assign p[13][26] = x[13]&y[13];
assign p[13][27] = x[14]&y[13];
assign p[13][28] = x[15]&y[13];
assign p[13][29] = x[16]&y[13];
assign p[13][30] = x[17]&y[13];
assign p[13][31] = x[18]&y[13];
assign p[13][32] = x[19]&y[13];
assign p[13][33] = x[20]&y[13];
assign p[13][34] = x[21]&y[13];
assign p[13][35] = x[22]&y[13];
assign p[13][36] = x[23]&y[13];
assign p[13][37] = x[24]&y[13];
assign p[13][38] = x[25]&y[13];
assign p[13][39] = x[26]&y[13];
assign p[13][40] = x[27]&y[13];
assign p[13][41] = x[28]&y[13];
assign p[13][42] = x[29]&y[13];
assign p[13][43] = x[30]&y[13];
assign p[13][44] = x[31]&y[13];
assign p[13][63:45] =1'b0;

//level 15
assign p[14][13:0]= 1'b0;
assign p[14][14] = x[0] & y[14];
assign p[14][15] = x[1]&y[14];
assign p[14][16] = x[2]&y[14];
assign p[14][17] = x[3]&y[14];
assign p[14][18] = x[4]&y[14];
assign p[14][19] = x[5]&y[14];
assign p[14][20] = x[6]&y[14];
assign p[14][21] = x[7]&y[14];
assign p[14][22] = x[8]&y[14];
assign p[14][23] = x[9]&y[14];
assign p[14][24] = x[10]&y[14];
assign p[14][25] = x[11]&y[14];
assign p[14][26] = x[12]&y[14];
assign p[14][27] = x[13]&y[14];
assign p[14][28] = x[14]&y[14];
assign p[14][29] = x[15]&y[14];
assign p[14][30] = x[16]&y[14];
assign p[14][31] = x[17]&y[14];
assign p[14][32] = x[18]&y[14];
assign p[14][33] = x[19]&y[14];
assign p[14][34] = x[20]&y[14];
assign p[14][35] = x[21]&y[14];
assign p[14][36] = x[22]&y[14];
assign p[14][37] = x[23]&y[14];
assign p[14][38] = x[24]&y[14];
assign p[14][39] = x[25]&y[14];
assign p[14][40] = x[26]&y[14];
assign p[14][41] = x[27]&y[14];
assign p[14][42] = x[28]&y[14];
assign p[14][43] = x[29]&y[14];
assign p[14][44] = x[30]&y[14];
assign p[14][45] = x[31]&y[14];
assign p[14][63:46] =1'b0;

//level 16
assign p[15][14:0]= 1'b0;
assign p[15][15] = x[0] & y[15];
assign p[15][16] = x[1]&y[15];
assign p[15][17] = x[2]&y[15];
assign p[15][18] = x[3]&y[15];
assign p[15][19] = x[4]&y[15];
assign p[15][20] = x[5]&y[15];
assign p[15][21] = x[6]&y[15];
assign p[15][22] = x[7]&y[15];
assign p[15][23] = x[8]&y[15];
assign p[15][24] = x[9]&y[15];
assign p[15][25] = x[10]&y[15];
assign p[15][26] = x[11]&y[15];
assign p[15][27] = x[12]&y[15];
assign p[15][28] = x[13]&y[15];
assign p[15][29] = x[14]&y[15];
assign p[15][30] = x[15]&y[15];
assign p[15][31] = x[16]&y[15];
assign p[15][32] = x[17]&y[15];
assign p[15][33] = x[18]&y[15];
assign p[15][34] = x[19]&y[15];
assign p[15][35] = x[20]&y[15];
assign p[15][36] = x[21]&y[15];
assign p[15][37] = x[22]&y[15];
assign p[15][38] = x[23]&y[15];
assign p[15][39] = x[24]&y[15];
assign p[15][40] = x[25]&y[15];
assign p[15][41] = x[26]&y[15];
assign p[15][42] = x[27]&y[15];
assign p[15][43] = x[28]&y[15];
assign p[15][44] = x[29]&y[15];
assign p[15][45] = x[30]&y[15];
assign p[15][46] = x[31]&y[15];
assign p[15][63:47] =1'b0;

//level 17
assign p[16][15:0]= 1'b0;
assign p[16][16] = x[0] & y[16];
assign p[16][17] = x[1]&y[16];
assign p[16][18] = x[2]&y[16];
assign p[16][19] = x[3]&y[16];
assign p[16][20] = x[4]&y[16];
assign p[16][21] = x[5]&y[16];
assign p[16][22] = x[6]&y[16];
assign p[16][23] = x[7]&y[16];
assign p[16][24] = x[8]&y[16];
assign p[16][25] = x[9]&y[16];
assign p[16][26] = x[10]&y[16];
assign p[16][27] = x[11]&y[16];
assign p[16][28] = x[12]&y[16];
assign p[16][29] = x[13]&y[16];
assign p[16][30] = x[14]&y[16];
assign p[16][31] = x[15]&y[16];
assign p[16][32] = x[16]&y[16];
assign p[16][33] = x[17]&y[16];
assign p[16][34] = x[18]&y[16];
assign p[16][35] = x[19]&y[16];
assign p[16][36] = x[20]&y[16];
assign p[16][37] = x[21]&y[16];
assign p[16][38] = x[22]&y[16];
assign p[16][39] = x[23]&y[16];
assign p[16][40] = x[24]&y[16];
assign p[16][41] = x[25]&y[16];
assign p[16][42] = x[26]&y[16];
assign p[16][43] = x[27]&y[16];
assign p[16][44] = x[28]&y[16];
assign p[16][45] = x[29]&y[16];
assign p[16][46] = x[30]&y[16];
assign p[16][47] = x[31]&y[16];
assign p[16][63:48] =1'b0;

//level 18
assign p[17][16:0]= 1'b0;
assign p[17][17] = x[0] & y[17];
assign p[17][18] = x[1]&y[17];
assign p[17][19] = x[2]&y[17];
assign p[17][20] = x[3]&y[17];
assign p[17][21] = x[4]&y[17];
assign p[17][22] = x[5]&y[17];
assign p[17][23] = x[6]&y[17];
assign p[17][24] = x[7]&y[17];
assign p[17][25] = x[8]&y[17];
assign p[17][26] = x[9]&y[17];
assign p[17][27] = x[10]&y[17];
assign p[17][28] = x[11]&y[17];
assign p[17][29] = x[12]&y[17];
assign p[17][30] = x[13]&y[17];
assign p[17][31] = x[14]&y[17];
assign p[17][32] = x[15]&y[17];
assign p[17][33] = x[16]&y[17];
assign p[17][34] = x[17]&y[17];
assign p[17][35] = x[18]&y[17];
assign p[17][36] = x[19]&y[17];
assign p[17][37] = x[20]&y[17];
assign p[17][38] = x[21]&y[17];
assign p[17][39] = x[22]&y[17];
assign p[17][40] = x[23]&y[17];
assign p[17][41] = x[24]&y[17];
assign p[17][42] = x[25]&y[17];
assign p[17][43] = x[26]&y[17];
assign p[17][44] = x[27]&y[17];
assign p[17][45] = x[28]&y[17];
assign p[17][46] = x[29]&y[17];
assign p[17][47] = x[30]&y[17];
assign p[17][48] = x[31]&y[17];
assign p[17][63:49] =1'b0;

//level 19
assign p[18][17:0]= 1'b0;
assign p[18][18] = x[0] & y[18];
assign p[18][19] = x[1]&y[18];
assign p[18][20] = x[2]&y[18];
assign p[18][21] = x[3]&y[18];
assign p[18][22] = x[4]&y[18];
assign p[18][23] = x[5]&y[18];
assign p[18][24] = x[6]&y[18];
assign p[18][25] = x[7]&y[18];
assign p[18][26] = x[8]&y[18];
assign p[18][27] = x[9]&y[18];
assign p[18][28] = x[10]&y[18];
assign p[18][29] = x[11]&y[18];
assign p[18][30] = x[12]&y[18];
assign p[18][31] = x[13]&y[18];
assign p[18][32] = x[14]&y[18];
assign p[18][33] = x[15]&y[18];
assign p[18][34] = x[16]&y[18];
assign p[18][35] = x[17]&y[18];
assign p[18][36] = x[18]&y[18];
assign p[18][37] = x[19]&y[18];
assign p[18][38] = x[20]&y[18];
assign p[18][39] = x[21]&y[18];
assign p[18][40] = x[22]&y[18];
assign p[18][41] = x[23]&y[18];
assign p[18][42] = x[24]&y[18];
assign p[18][43] = x[25]&y[18];
assign p[18][44] = x[26]&y[18];
assign p[18][45] = x[27]&y[18];
assign p[18][46] = x[28]&y[18];
assign p[18][47] = x[29]&y[18];
assign p[18][48] = x[30]&y[18];
assign p[18][49] = x[31]&y[18];
assign p[18][63:50] =1'b0;

//level 20
assign p[19][18:0]= 1'b0;
assign p[19][19] = x[0] & y[19];
assign p[19][20] = x[1]&y[19];
assign p[19][21] = x[2]&y[19];
assign p[19][22] = x[3]&y[19];
assign p[19][23] = x[4]&y[19];
assign p[19][24] = x[5]&y[19];
assign p[19][25] = x[6]&y[19];
assign p[19][26] = x[7]&y[19];
assign p[19][27] = x[8]&y[19];
assign p[19][28] = x[9]&y[19];
assign p[19][29] = x[10]&y[19];
assign p[19][30] = x[11]&y[19];
assign p[19][31] = x[12]&y[19];
assign p[19][32] = x[13]&y[19];
assign p[19][33] = x[14]&y[19];
assign p[19][34] = x[15]&y[19];
assign p[19][35] = x[16]&y[19];
assign p[19][36] = x[17]&y[19];
assign p[19][37] = x[18]&y[19];
assign p[19][38] = x[19]&y[19];
assign p[19][39] = x[20]&y[19];
assign p[19][40] = x[21]&y[19];
assign p[19][41] = x[22]&y[19];
assign p[19][42] = x[23]&y[19];
assign p[19][43] = x[24]&y[19];
assign p[19][44] = x[25]&y[19];
assign p[19][45] = x[26]&y[19];
assign p[19][46] = x[27]&y[19];
assign p[19][47] = x[28]&y[19];
assign p[19][48] = x[29]&y[19];
assign p[19][49] = x[30]&y[19];
assign p[19][50] = x[31]&y[19];
assign p[19][63:51] =1'b0;

//level 21
assign p[20][19:0]= 1'b0;
assign p[20][20] = x[0] & y[20];
assign p[20][21] = x[1]&y[20];
assign p[20][22] = x[2]&y[20];
assign p[20][23] = x[3]&y[20];
assign p[20][24] = x[4]&y[20];
assign p[20][25] = x[5]&y[20];
assign p[20][26] = x[6]&y[20];
assign p[20][27] = x[7]&y[20];
assign p[20][28] = x[8]&y[20];
assign p[20][29] = x[9]&y[20];
assign p[20][30] = x[10]&y[20];
assign p[20][31] = x[11]&y[20];
assign p[20][32] = x[12]&y[20];
assign p[20][33] = x[13]&y[20];
assign p[20][34] = x[14]&y[20];
assign p[20][35] = x[15]&y[20];
assign p[20][36] = x[16]&y[20];
assign p[20][37] = x[17]&y[20];
assign p[20][38] = x[18]&y[20];
assign p[20][39] = x[19]&y[20];
assign p[20][40] = x[20]&y[20];
assign p[20][41] = x[21]&y[20];
assign p[20][42] = x[22]&y[20];
assign p[20][43] = x[23]&y[20];
assign p[20][44] = x[24]&y[20];
assign p[20][45] = x[25]&y[20];
assign p[20][46] = x[26]&y[20];
assign p[20][47] = x[27]&y[20];
assign p[20][48] = x[28]&y[20];
assign p[20][49] = x[29]&y[20];
assign p[20][50] = x[30]&y[20];
assign p[20][51] = x[31]&y[20];
assign p[20][63:52] =1'b0;

//level 22
assign p[21][20:0]= 1'b0;
assign p[21][21] = x[0] & y[21];
assign p[21][22] = x[1]&y[21];
assign p[21][23] = x[2]&y[21];
assign p[21][24] = x[3]&y[21];
assign p[21][25] = x[4]&y[21];
assign p[21][26] = x[5]&y[21];
assign p[21][27] = x[6]&y[21];
assign p[21][28] = x[7]&y[21];
assign p[21][29] = x[8]&y[21];
assign p[21][30] = x[9]&y[21];
assign p[21][31] = x[10]&y[21];
assign p[21][32] = x[11]&y[21];
assign p[21][33] = x[12]&y[21];
assign p[21][34] = x[13]&y[21];
assign p[21][35] = x[14]&y[21];
assign p[21][36] = x[15]&y[21];
assign p[21][37] = x[16]&y[21];
assign p[21][38] = x[17]&y[21];
assign p[21][39] = x[18]&y[21];
assign p[21][40] = x[19]&y[21];
assign p[21][41] = x[20]&y[21];
assign p[21][42] = x[21]&y[21];
assign p[21][43] = x[22]&y[21];
assign p[21][44] = x[23]&y[21];
assign p[21][45] = x[24]&y[21];
assign p[21][46] = x[25]&y[21];
assign p[21][47] = x[26]&y[21];
assign p[21][48] = x[27]&y[21];
assign p[21][49] = x[28]&y[21];
assign p[21][50] = x[29]&y[21];
assign p[21][51] = x[30]&y[21];
assign p[21][52] = x[31]&y[21];
assign p[21][63:53] =1'b0;

//level 23
assign p[22][21:0]= 1'b0;
assign p[22][22] = x[0] & y[22];
assign p[22][23] = x[1]&y[22];
assign p[22][24] = x[2]&y[22];
assign p[22][25] = x[3]&y[22];
assign p[22][26] = x[4]&y[22];
assign p[22][27] = x[5]&y[22];
assign p[22][28] = x[6]&y[22];
assign p[22][29] = x[7]&y[22];
assign p[22][30] = x[8]&y[22];
assign p[22][31] = x[9]&y[22];
assign p[22][32] = x[10]&y[22];
assign p[22][33] = x[11]&y[22];
assign p[22][34] = x[12]&y[22];
assign p[22][35] = x[13]&y[22];
assign p[22][36] = x[14]&y[22];
assign p[22][37] = x[15]&y[22];
assign p[22][38] = x[16]&y[22];
assign p[22][39] = x[17]&y[22];
assign p[22][40] = x[18]&y[22];
assign p[22][41] = x[19]&y[22];
assign p[22][42] = x[20]&y[22];
assign p[22][43] = x[21]&y[22];
assign p[22][44] = x[22]&y[22];
assign p[22][45] = x[23]&y[22];
assign p[22][46] = x[24]&y[22];
assign p[22][47] = x[25]&y[22];
assign p[22][48] = x[26]&y[22];
assign p[22][49] = x[27]&y[22];
assign p[22][50] = x[28]&y[22];
assign p[22][51] = x[29]&y[22];
assign p[22][52] = x[30]&y[22];
assign p[22][53] = x[31]&y[22];
assign p[22][63:54] =1'b0;

//level 24
assign p[23][22:0]= 1'b0;
assign p[23][23] = x[0] & y[23];
assign p[23][24] = x[1]&y[23];
assign p[23][25] = x[2]&y[23];
assign p[23][26] = x[3]&y[23];
assign p[23][27] = x[4]&y[23];
assign p[23][28] = x[5]&y[23];
assign p[23][29] = x[6]&y[23];
assign p[23][30] = x[7]&y[23];
assign p[23][31] = x[8]&y[23];
assign p[23][32] = x[9]&y[23];
assign p[23][33] = x[10]&y[23];
assign p[23][34] = x[11]&y[23];
assign p[23][35] = x[12]&y[23];
assign p[23][36] = x[13]&y[23];
assign p[23][37] = x[14]&y[23];
assign p[23][38] = x[15]&y[23];
assign p[23][39] = x[16]&y[23];
assign p[23][40] = x[17]&y[23];
assign p[23][41] = x[18]&y[23];
assign p[23][42] = x[19]&y[23];
assign p[23][43] = x[20]&y[23];
assign p[23][44] = x[21]&y[23];
assign p[23][45] = x[22]&y[23];
assign p[23][46] = x[23]&y[23];
assign p[23][47] = x[24]&y[23];
assign p[23][48] = x[25]&y[23];
assign p[23][49] = x[26]&y[23];
assign p[23][50] = x[27]&y[23];
assign p[23][51] = x[28]&y[23];
assign p[23][52] = x[29]&y[23];
assign p[23][53] = x[30]&y[23];
assign p[23][54] = x[31]&y[23];
assign p[23][63:55] =1'b0;

//level 25
assign p[24][23:0]= 1'b0;
assign p[24][24] = x[0] & y[24];
assign p[24][25] = x[1]&y[24];
assign p[24][26] = x[2]&y[24];
assign p[24][27] = x[3]&y[24];
assign p[24][28] = x[4]&y[24];
assign p[24][29] = x[5]&y[24];
assign p[24][30] = x[6]&y[24];
assign p[24][31] = x[7]&y[24];
assign p[24][32] = x[8]&y[24];
assign p[24][33] = x[9]&y[24];
assign p[24][34] = x[10]&y[24];
assign p[24][35] = x[11]&y[24];
assign p[24][36] = x[12]&y[24];
assign p[24][37] = x[13]&y[24];
assign p[24][38] = x[14]&y[24];
assign p[24][39] = x[15]&y[24];
assign p[24][40] = x[16]&y[24];
assign p[24][41] = x[17]&y[24];
assign p[24][42] = x[18]&y[24];
assign p[24][43] = x[19]&y[24];
assign p[24][44] = x[20]&y[24];
assign p[24][45] = x[21]&y[24];
assign p[24][46] = x[22]&y[24];
assign p[24][47] = x[23]&y[24];
assign p[24][48] = x[24]&y[24];
assign p[24][49] = x[25]&y[24];
assign p[24][50] = x[26]&y[24];
assign p[24][51] = x[27]&y[24];
assign p[24][52] = x[28]&y[24];
assign p[24][53] = x[29]&y[24];
assign p[24][54] = x[30]&y[24];
assign p[24][55] = x[31]&y[24];
assign p[24][63:56] =1'b0;

//level 26
assign p[25][24:0]= 1'b0;
assign p[25][25] = x[0] & y[25];
assign p[25][26] = x[1]&y[25];
assign p[25][27] = x[2]&y[25];
assign p[25][28] = x[3]&y[25];
assign p[25][29] = x[4]&y[25];
assign p[25][30] = x[5]&y[25];
assign p[25][31] = x[6]&y[25];
assign p[25][32] = x[7]&y[25];
assign p[25][33] = x[8]&y[25];
assign p[25][34] = x[9]&y[25];
assign p[25][35] = x[10]&y[25];
assign p[25][36] = x[11]&y[25];
assign p[25][37] = x[12]&y[25];
assign p[25][38] = x[13]&y[25];
assign p[25][39] = x[14]&y[25];
assign p[25][40] = x[15]&y[25];
assign p[25][41] = x[16]&y[25];
assign p[25][42] = x[17]&y[25];
assign p[25][43] = x[18]&y[25];
assign p[25][44] = x[19]&y[25];
assign p[25][45] = x[20]&y[25];
assign p[25][46] = x[21]&y[25];
assign p[25][47] = x[22]&y[25];
assign p[25][48] = x[23]&y[25];
assign p[25][49] = x[24]&y[25];
assign p[25][50] = x[25]&y[25];
assign p[25][51] = x[26]&y[25];
assign p[25][52] = x[27]&y[25];
assign p[25][53] = x[28]&y[25];
assign p[25][54] = x[29]&y[25];
assign p[25][55] = x[30]&y[25];
assign p[25][56] = x[31]&y[25];
assign p[25][63:57] =1'b0;

//level 27
assign p[26][25:0]= 1'b0;
assign p[26][26] = x[0] & y[26];
assign p[26][27] = x[1]&y[26];
assign p[26][28] = x[2]&y[26];
assign p[26][29] = x[3]&y[26];
assign p[26][30] = x[4]&y[26];
assign p[26][31] = x[5]&y[26];
assign p[26][32] = x[6]&y[26];
assign p[26][33] = x[7]&y[26];
assign p[26][34] = x[8]&y[26];
assign p[26][35] = x[9]&y[26];
assign p[26][36] = x[10]&y[26];
assign p[26][37] = x[11]&y[26];
assign p[26][38] = x[12]&y[26];
assign p[26][39] = x[13]&y[26];
assign p[26][40] = x[14]&y[26];
assign p[26][41] = x[15]&y[26];
assign p[26][42] = x[16]&y[26];
assign p[26][43] = x[17]&y[26];
assign p[26][44] = x[18]&y[26];
assign p[26][45] = x[19]&y[26];
assign p[26][46] = x[20]&y[26];
assign p[26][47] = x[21]&y[26];
assign p[26][48] = x[22]&y[26];
assign p[26][49] = x[23]&y[26];
assign p[26][50] = x[24]&y[26];
assign p[26][51] = x[25]&y[26];
assign p[26][52] = x[26]&y[26];
assign p[26][53] = x[27]&y[26];
assign p[26][54] = x[28]&y[26];
assign p[26][55] = x[29]&y[26];
assign p[26][56] = x[30]&y[26];
assign p[26][57] = x[31]&y[26];
assign p[26][63:58] =1'b0;

//level 28
assign p[27][26:0]= 1'b0;
assign p[27][27] = x[0] & y[27];
assign p[27][28] = x[1]&y[27];
assign p[27][29] = x[2]&y[27];
assign p[27][30] = x[3]&y[27];
assign p[27][31] = x[4]&y[27];
assign p[27][32] = x[5]&y[27];
assign p[27][33] = x[6]&y[27];
assign p[27][34] = x[7]&y[27];
assign p[27][35] = x[8]&y[27];
assign p[27][36] = x[9]&y[27];
assign p[27][37] = x[10]&y[27];
assign p[27][38] = x[11]&y[27];
assign p[27][39] = x[12]&y[27];
assign p[27][40] = x[13]&y[27];
assign p[27][41] = x[14]&y[27];
assign p[27][42] = x[15]&y[27];
assign p[27][43] = x[16]&y[27];
assign p[27][44] = x[17]&y[27];
assign p[27][45] = x[18]&y[27];
assign p[27][46] = x[19]&y[27];
assign p[27][47] = x[20]&y[27];
assign p[27][48] = x[21]&y[27];
assign p[27][49] = x[22]&y[27];
assign p[27][50] = x[23]&y[27];
assign p[27][51] = x[24]&y[27];
assign p[27][52] = x[25]&y[27];
assign p[27][53] = x[26]&y[27];
assign p[27][54] = x[27]&y[27];
assign p[27][55] = x[28]&y[27];
assign p[27][56] = x[29]&y[27];
assign p[27][57] = x[30]&y[27];
assign p[27][58] = x[31]&y[27];
assign p[27][63:59] =1'b0;

//level 29
assign p[28][27:0]= 1'b0;
assign p[28][28] = x[0] & y[28];
assign p[28][29] = x[1]&y[28];
assign p[28][30] = x[2]&y[28];
assign p[28][31] = x[3]&y[28];
assign p[28][32] = x[4]&y[28];
assign p[28][33] = x[5]&y[28];
assign p[28][34] = x[6]&y[28];
assign p[28][35] = x[7]&y[28];
assign p[28][36] = x[8]&y[28];
assign p[28][37] = x[9]&y[28];
assign p[28][38] = x[10]&y[28];
assign p[28][39] = x[11]&y[28];
assign p[28][40] = x[12]&y[28];
assign p[28][41] = x[13]&y[28];
assign p[28][42] = x[14]&y[28];
assign p[28][43] = x[15]&y[28];
assign p[28][44] = x[16]&y[28];
assign p[28][45] = x[17]&y[28];
assign p[28][46] = x[18]&y[28];
assign p[28][47] = x[19]&y[28];
assign p[28][48] = x[20]&y[28];
assign p[28][49] = x[21]&y[28];
assign p[28][50] = x[22]&y[28];
assign p[28][51] = x[23]&y[28];
assign p[28][52] = x[24]&y[28];
assign p[28][53] = x[25]&y[28];
assign p[28][54] = x[26]&y[28];
assign p[28][55] = x[27]&y[28];
assign p[28][56] = x[28]&y[28];
assign p[28][57] = x[29]&y[28];
assign p[28][58] = x[30]&y[28];
assign p[28][59] = x[31]&y[28];
assign p[28][63:60] =1'b0;

//level 30
assign p[29][28:0]= 1'b0;
assign p[29][29] = x[0] & y[29];
assign p[29][30] = x[1]&y[29];
assign p[29][31] = x[2]&y[29];
assign p[29][32] = x[3]&y[29];
assign p[29][33] = x[4]&y[29];
assign p[29][34] = x[5]&y[29];
assign p[29][35] = x[6]&y[29];
assign p[29][36] = x[7]&y[29];
assign p[29][37] = x[8]&y[29];
assign p[29][38] = x[9]&y[29];
assign p[29][39] = x[10]&y[29];
assign p[29][40] = x[11]&y[29];
assign p[29][41] = x[12]&y[29];
assign p[29][42] = x[13]&y[29];
assign p[29][43] = x[14]&y[29];
assign p[29][44] = x[15]&y[29];
assign p[29][45] = x[16]&y[29];
assign p[29][46] = x[17]&y[29];
assign p[29][47] = x[18]&y[29];
assign p[29][48] = x[19]&y[29];
assign p[29][49] = x[20]&y[29];
assign p[29][50] = x[21]&y[29];
assign p[29][51] = x[22]&y[29];
assign p[29][52] = x[23]&y[29];
assign p[29][53] = x[24]&y[29];
assign p[29][54] = x[25]&y[29];
assign p[29][55] = x[26]&y[29];
assign p[29][56] = x[27]&y[29];
assign p[29][57] = x[28]&y[29];
assign p[29][58] = x[29]&y[29];
assign p[29][59] = x[30]&y[29];
assign p[29][60] = x[31]&y[29];
assign p[29][63:61] =1'b0;

//level 31
assign p[30][29:0]= 1'b0;
assign p[30][30] = x[0] & y[30];
assign p[30][31] = x[1]&y[30];
assign p[30][32] = x[2]&y[30];
assign p[30][33] = x[3]&y[30];
assign p[30][34] = x[4]&y[30];
assign p[30][35] = x[5]&y[30];
assign p[30][36] = x[6]&y[30];
assign p[30][37] = x[7]&y[30];
assign p[30][38] = x[8]&y[30];
assign p[30][39] = x[9]&y[30];
assign p[30][40] = x[10]&y[30];
assign p[30][41] = x[11]&y[30];
assign p[30][42] = x[12]&y[30];
assign p[30][43] = x[13]&y[30];
assign p[30][44] = x[14]&y[30];
assign p[30][45] = x[15]&y[30];
assign p[30][46] = x[16]&y[30];
assign p[30][47] = x[17]&y[30];
assign p[30][48] = x[18]&y[30];
assign p[30][49] = x[19]&y[30];
assign p[30][50] = x[20]&y[30];
assign p[30][51] = x[21]&y[30];
assign p[30][52] = x[22]&y[30];
assign p[30][53] = x[23]&y[30];
assign p[30][54] = x[24]&y[30];
assign p[30][55] = x[25]&y[30];
assign p[30][56] = x[26]&y[30];
assign p[30][57] = x[27]&y[30];
assign p[30][58] = x[28]&y[30];
assign p[30][59] = x[29]&y[30];
assign p[30][60] = x[30]&y[30];
assign p[30][61] = x[31]&y[30];
assign p[30][63:62] =1'b0;

//level 32
assign p[31][30:0]= 1'b0;
assign p[31][31] = x[0] & y[31];
assign p[31][32] = x[1]&y[31];
assign p[31][33] = x[2]&y[31];
assign p[31][34] = x[3]&y[31];
assign p[31][35] = x[4]&y[31];
assign p[31][36] = x[5]&y[31];
assign p[31][37] = x[6]&y[31];
assign p[31][38] = x[7]&y[31];
assign p[31][39] = x[8]&y[31];
assign p[31][40] = x[9]&y[31];
assign p[31][41] = x[10]&y[31];
assign p[31][42] = x[11]&y[31];
assign p[31][43] = x[12]&y[31];
assign p[31][44] = x[13]&y[31];
assign p[31][45] = x[14]&y[31];
assign p[31][46] = x[15]&y[31];
assign p[31][47] = x[16]&y[31];
assign p[31][48] = x[17]&y[31];
assign p[31][49] = x[18]&y[31];
assign p[31][50] = x[19]&y[31];
assign p[31][51] = x[20]&y[31];
assign p[31][52] = x[21]&y[31];
assign p[31][53] = x[22]&y[31];
assign p[31][54] = x[23]&y[31];
assign p[31][55] = x[24]&y[31];
assign p[31][56] = x[25]&y[31];
assign p[31][57] = x[26]&y[31];
assign p[31][58] = x[27]&y[31];
assign p[31][59] = x[28]&y[31];
assign p[31][60] = x[29]&y[31];
assign p[31][61] = x[30]&y[31];
assign p[31][62] = x[31]&y[31];
assign p[31][63] = 1'b0;

//Stage1(32/3 ~ 10)
csa a1(p[0],p[1],p[2],s1,c1);
csa a2(p[3],p[4],p[5],s2,c2);
csa a3(p[6],p[7],p[8],s3,c3);
csa a4(p[9],p[10],p[11],s4,c4);
csa a5(p[12],p[13],p[14],s5,c5);
csa a6(p[15],p[16],p[17],s6,c6);
csa a7(p[18],p[19],p[20],s7,c7);
csa a8(p[21],p[22],p[23],s8,c8);
csa a9(p[24],p[25],p[26],s9,c9);
csa a10(p[27],p[28],p[29],s10,c10);
//csa a11(p[30],p[31],64'd0,c10[64],s11,c11);

//Stage2(20/3 ~ 7)
csa a11(s1,c1,s2,s11,c11);
csa a12(c2,s3,c3,s12,c12);
csa a13(s4,c4,s5,s13,c13);
csa a14(c5,s6,c6,s14,c14);
csa a15(s7,c7,s8,s15,c15);
csa a16(c8,s9,c9,s16,c16);
csa a17(s10,c10,p[30],s17,c17);

//Stage3(14/3 ~ 5)
csa a18(s11,c11,s12,s18,c18);
csa a19(c12,s13,c13,s19,c19);
csa a20(s14,c14,s15,s20,c20);
csa a21(c15,s16,c16,s21,c21);
csa a22(s17,c17,p[31],s22,c22);

//Stage4(10/3 ~3)
csa a23(s18,c18,s19,s23,c23);
csa a24(c19,s20,c20,s24,c24);
csa a25(s21,c21,s22,s25,c25);

//Stage5(6/3 ~2)
csa a26(c22,s23,c23,s26,c26);
csa a27(s24,c24,s25,s27,c27);

//Stage6(4/3 ~1)
csa a28(c25,s26,c26,s28,c28);

csa a29(s27,c27,s28,s29,c29);

csa a30(c28,s29,c29,s30,c30);

pre32 p1(o[31:0],cout1,s30[31:0],c30[31:0],1'b0);
pre32 p2(o[63:32],cout2,s30[63:32],c30[63:32],cout1);

assign o[64]=cout2;
endmodule