module multiplier_tb();

reg [31:0]num1,num2;
wire [31:0]num3;
/*//sign bit
reg s1,s2;
wire s3;
//exponent
reg [7:0]exp1,exp2;
wire [7:0]exp3;
//mantissa
reg [22:0]man1,man2;
wire [22:0]man3;
reg [22:0]m1,m2;*/

fpmultiplier m(num1,num2,num3);

initial 
begin
num1=32'b11000001100101000000000000000000;
num2=32'b01000001000110000000000000000000;

//num1=32'd12;
//num2=32'd3;
//9.5
// 1  10000110  01011111100000000000000  //-175.75
#5
num1=32'b10111111110000000000000000000000;       
num2=32'b10111111110000000000000000000000;
//-1.5          
// 0  10000000  00100000000000000000000
#5                                     
num1=32'b00111111110000000000000000000000; 
num1=32'b11000001000110000000000000000000;       
//-9.5                                   
// 0  10000010  11001000000000000000000  
#5
num1=32'b11000001100101000000000000000000;
//-18.5
num2=32'b11000011101010110010000000000000;
#5
num1=32'b01111111111111111111111111111111;
num2=32'b01111111111111111111111111111111;
#5
num1=32'b01000111110110110101110010010000;
num2=32'b01000111110110110101110010010000;
#5
num1=32'b01000111110110110101110010010000;
num2=32'b11001000000000010101010010010000;
end

initial
begin
$monitor($time,"  num1=%b,\n\t\t      num2=%b,\n\t\t      num3=%b",num1,num2,num3);
end
endmodule