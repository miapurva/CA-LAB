//`include "../FPM/FPM.v"

module FPM_TB();

	reg[31:0] A,B;
	reg clk;

	wire[31:0] SUM;

	FPM float_mult(A,B,SUM,clk);

	always #2 clk=~clk;

	initial
	begin
		clk=0;

		#1 A=32'b11000001100100000000000000000000;
		   B=32'b01000001000110000000000000000000;

		 #4 A=32'b01000010111101110000000000000000;
		 	B=32'b11000001010010000000000000000000;

		 #4 A=32'b00111111101000000000000000000000; //1.25
		 	B=32'b00111110100110011001100110011001; //0.3

		 #4 A=32'b01000100011110100000000000000000; //1000
		 	B=32'b00111111000000000000000000000000; //0.5

		 #4 A=32'b01000100011110100000000000000000; //1000
		 	B=32'b00111110010011001100110011001100; //0.2

		 #4 A=32'b11000001001000111100000010100100; //10.234532121
		 	B=32'b01000100011111111101110100000001; //1023.4532121

		 #4 A=32'b00111111000000000000000000000000; //0.5
		 	B=32'b00110111001001111100010110101100; //0.00001

		#100 $finish;
	end

	initial
	begin
		$monitor($time," A=%b B=%b SUM=%h",A,B,SUM);
	end
endmodule // FPM